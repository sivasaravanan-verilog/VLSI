
typedef class karthik;
  
  class kaviya;
    karthik k;
  endclass
  
  class karthik;
    kaviya v;
  endclass
  
  
  module love;
    
    initial begin
      karthik c1;
      kaviya v1;
      
      $display("*******************");
      $display("\n typedef class");
      $display("\n remove compiler error");
    end
  endmodule
