interface inter;
  logic clk;
  logic rst;
  logic [7:0] data;
  logic [7:0] dout;
  logic wen,ren;
  logic full, empty;
endinterface
