module andg (A, B, Y); 
  input A,B; 
  output Y; 
  and(A,B);
endmodule
