class transaction;
  bit clk;
  bit[8:0]wdata;
  bit[8:0]addr;
  bit wen;
  bit[8:0]rdata;
endclass
