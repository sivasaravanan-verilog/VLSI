interface i2c_interface() ;
	logic scl_pad_i ;   
	logic scl_pad_o  ;  
	logic scl_padoen_o ;
	logic sda_pad_i   ;
	logic sda_pad_o   ;
	logic sda_padoen_o ;

endinterface
