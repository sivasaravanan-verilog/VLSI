module simple_function();
  
   function  myfunction;
   input a, b, c, d;
   begin
     myfunction = ((a+b) + (c-d));
   end
   endfunction
   
  endmodule
