module org(A,B,Y); 
  input A,B; 
  output Y; 
  or(Y,A,B);
endmodule
