import uvm_pkg::*;
`include "uvm_macros.svh"

`include "apb_2_i2c_defines.sv"
`include "apb_transaction.sv"
`include "apb_sequence.sv"
`include "apb_sequencer.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_agent.sv"

`include "i2c_transaction.sv"
`include "i2c_monitor.sv"
`include "i2c_agent.sv"
`include "apb_2_i2c_sb.sv"
`include "apb_2_i2c_env.sv"
`include "apb_2_i2c_test.sv"

